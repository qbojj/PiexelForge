// HPS.v

// Generated using ACDS version 24.1 1077

`timescale 1 ps / 1 ps
module HPS (
		input  wire        f2h_sdram_clk_clk,       //   f2h_sdram_clk.clk
		input  wire [31:0] f2h_sdram_slave_araddr,  // f2h_sdram_slave.araddr
		input  wire [3:0]  f2h_sdram_slave_arlen,   //                .arlen
		input  wire [7:0]  f2h_sdram_slave_arid,    //                .arid
		input  wire [2:0]  f2h_sdram_slave_arsize,  //                .arsize
		input  wire [1:0]  f2h_sdram_slave_arburst, //                .arburst
		input  wire [1:0]  f2h_sdram_slave_arlock,  //                .arlock
		input  wire [2:0]  f2h_sdram_slave_arprot,  //                .arprot
		input  wire        f2h_sdram_slave_arvalid, //                .arvalid
		input  wire [3:0]  f2h_sdram_slave_arcache, //                .arcache
		input  wire [31:0] f2h_sdram_slave_awaddr,  //                .awaddr
		input  wire [3:0]  f2h_sdram_slave_awlen,   //                .awlen
		input  wire [7:0]  f2h_sdram_slave_awid,    //                .awid
		input  wire [2:0]  f2h_sdram_slave_awsize,  //                .awsize
		input  wire [1:0]  f2h_sdram_slave_awburst, //                .awburst
		input  wire [1:0]  f2h_sdram_slave_awlock,  //                .awlock
		input  wire [2:0]  f2h_sdram_slave_awprot,  //                .awprot
		input  wire        f2h_sdram_slave_awvalid, //                .awvalid
		input  wire [3:0]  f2h_sdram_slave_awcache, //                .awcache
		output wire [1:0]  f2h_sdram_slave_bresp,   //                .bresp
		output wire [7:0]  f2h_sdram_slave_bid,     //                .bid
		output wire        f2h_sdram_slave_bvalid,  //                .bvalid
		input  wire        f2h_sdram_slave_bready,  //                .bready
		output wire        f2h_sdram_slave_arready, //                .arready
		output wire        f2h_sdram_slave_awready, //                .awready
		input  wire        f2h_sdram_slave_rready,  //                .rready
		output wire [63:0] f2h_sdram_slave_rdata,   //                .rdata
		output wire [1:0]  f2h_sdram_slave_rresp,   //                .rresp
		output wire        f2h_sdram_slave_rlast,   //                .rlast
		output wire [7:0]  f2h_sdram_slave_rid,     //                .rid
		output wire        f2h_sdram_slave_rvalid,  //                .rvalid
		input  wire        f2h_sdram_slave_wlast,   //                .wlast
		input  wire        f2h_sdram_slave_wvalid,  //                .wvalid
		input  wire [63:0] f2h_sdram_slave_wdata,   //                .wdata
		input  wire [7:0]  f2h_sdram_slave_wstrb,   //                .wstrb
		output wire        f2h_sdram_slave_wready,  //                .wready
		input  wire [7:0]  f2h_sdram_slave_wid,     //                .wid
		input  wire        h2f_axi_clk_clk,         //     h2f_axi_clk.clk
		output wire [11:0] h2f_axi_master_awid,     //  h2f_axi_master.awid
		output wire [29:0] h2f_axi_master_awaddr,   //                .awaddr
		output wire [3:0]  h2f_axi_master_awlen,    //                .awlen
		output wire [2:0]  h2f_axi_master_awsize,   //                .awsize
		output wire [1:0]  h2f_axi_master_awburst,  //                .awburst
		output wire [1:0]  h2f_axi_master_awlock,   //                .awlock
		output wire [3:0]  h2f_axi_master_awcache,  //                .awcache
		output wire [2:0]  h2f_axi_master_awprot,   //                .awprot
		output wire        h2f_axi_master_awvalid,  //                .awvalid
		input  wire        h2f_axi_master_awready,  //                .awready
		output wire [11:0] h2f_axi_master_wid,      //                .wid
		output wire [31:0] h2f_axi_master_wdata,    //                .wdata
		output wire [3:0]  h2f_axi_master_wstrb,    //                .wstrb
		output wire        h2f_axi_master_wlast,    //                .wlast
		output wire        h2f_axi_master_wvalid,   //                .wvalid
		input  wire        h2f_axi_master_wready,   //                .wready
		input  wire [11:0] h2f_axi_master_bid,      //                .bid
		input  wire [1:0]  h2f_axi_master_bresp,    //                .bresp
		input  wire        h2f_axi_master_bvalid,   //                .bvalid
		output wire        h2f_axi_master_bready,   //                .bready
		output wire [11:0] h2f_axi_master_arid,     //                .arid
		output wire [29:0] h2f_axi_master_araddr,   //                .araddr
		output wire [3:0]  h2f_axi_master_arlen,    //                .arlen
		output wire [2:0]  h2f_axi_master_arsize,   //                .arsize
		output wire [1:0]  h2f_axi_master_arburst,  //                .arburst
		output wire [1:0]  h2f_axi_master_arlock,   //                .arlock
		output wire [3:0]  h2f_axi_master_arcache,  //                .arcache
		output wire [2:0]  h2f_axi_master_arprot,   //                .arprot
		output wire        h2f_axi_master_arvalid,  //                .arvalid
		input  wire        h2f_axi_master_arready,  //                .arready
		input  wire [11:0] h2f_axi_master_rid,      //                .rid
		input  wire [31:0] h2f_axi_master_rdata,    //                .rdata
		input  wire [1:0]  h2f_axi_master_rresp,    //                .rresp
		input  wire        h2f_axi_master_rlast,    //                .rlast
		input  wire        h2f_axi_master_rvalid,   //                .rvalid
		output wire        h2f_axi_master_rready,   //                .rready
		output wire        h2f_rst_reset_n,         //         h2f_rst.reset_n
		input  wire [31:0] irq0_irq,                //            irq0.irq
		input  wire [31:0] irq1_irq,                //            irq1.irq
		output wire [12:0] memory_mem_a,            //          memory.mem_a
		output wire [2:0]  memory_mem_ba,           //                .mem_ba
		output wire        memory_mem_ck,           //                .mem_ck
		output wire        memory_mem_ck_n,         //                .mem_ck_n
		output wire        memory_mem_cke,          //                .mem_cke
		output wire        memory_mem_cs_n,         //                .mem_cs_n
		output wire        memory_mem_ras_n,        //                .mem_ras_n
		output wire        memory_mem_cas_n,        //                .mem_cas_n
		output wire        memory_mem_we_n,         //                .mem_we_n
		output wire        memory_mem_reset_n,      //                .mem_reset_n
		inout  wire [31:0] memory_mem_dq,           //                .mem_dq
		inout  wire [3:0]  memory_mem_dqs,          //                .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,        //                .mem_dqs_n
		output wire        memory_mem_odt,          //                .mem_odt
		output wire [3:0]  memory_mem_dm,           //                .mem_dm
		input  wire        memory_oct_rzqin         //                .oct_rzqin
	);

	HPS_hps_0 #(
		.F2S_Width (0),
		.S2F_Width (1)
	) hps_0 (
		.mem_a              (memory_mem_a),            //           memory.mem_a
		.mem_ba             (memory_mem_ba),           //                 .mem_ba
		.mem_ck             (memory_mem_ck),           //                 .mem_ck
		.mem_ck_n           (memory_mem_ck_n),         //                 .mem_ck_n
		.mem_cke            (memory_mem_cke),          //                 .mem_cke
		.mem_cs_n           (memory_mem_cs_n),         //                 .mem_cs_n
		.mem_ras_n          (memory_mem_ras_n),        //                 .mem_ras_n
		.mem_cas_n          (memory_mem_cas_n),        //                 .mem_cas_n
		.mem_we_n           (memory_mem_we_n),         //                 .mem_we_n
		.mem_reset_n        (memory_mem_reset_n),      //                 .mem_reset_n
		.mem_dq             (memory_mem_dq),           //                 .mem_dq
		.mem_dqs            (memory_mem_dqs),          //                 .mem_dqs
		.mem_dqs_n          (memory_mem_dqs_n),        //                 .mem_dqs_n
		.mem_odt            (memory_mem_odt),          //                 .mem_odt
		.mem_dm             (memory_mem_dm),           //                 .mem_dm
		.oct_rzqin          (memory_oct_rzqin),        //                 .oct_rzqin
		.h2f_rst_n          (h2f_rst_reset_n),         //        h2f_reset.reset_n
		.f2h_sdram0_clk     (f2h_sdram_clk_clk),       // f2h_sdram0_clock.clk
		.f2h_sdram0_ARADDR  (f2h_sdram_slave_araddr),  //  f2h_sdram0_data.araddr
		.f2h_sdram0_ARLEN   (f2h_sdram_slave_arlen),   //                 .arlen
		.f2h_sdram0_ARID    (f2h_sdram_slave_arid),    //                 .arid
		.f2h_sdram0_ARSIZE  (f2h_sdram_slave_arsize),  //                 .arsize
		.f2h_sdram0_ARBURST (f2h_sdram_slave_arburst), //                 .arburst
		.f2h_sdram0_ARLOCK  (f2h_sdram_slave_arlock),  //                 .arlock
		.f2h_sdram0_ARPROT  (f2h_sdram_slave_arprot),  //                 .arprot
		.f2h_sdram0_ARVALID (f2h_sdram_slave_arvalid), //                 .arvalid
		.f2h_sdram0_ARCACHE (f2h_sdram_slave_arcache), //                 .arcache
		.f2h_sdram0_AWADDR  (f2h_sdram_slave_awaddr),  //                 .awaddr
		.f2h_sdram0_AWLEN   (f2h_sdram_slave_awlen),   //                 .awlen
		.f2h_sdram0_AWID    (f2h_sdram_slave_awid),    //                 .awid
		.f2h_sdram0_AWSIZE  (f2h_sdram_slave_awsize),  //                 .awsize
		.f2h_sdram0_AWBURST (f2h_sdram_slave_awburst), //                 .awburst
		.f2h_sdram0_AWLOCK  (f2h_sdram_slave_awlock),  //                 .awlock
		.f2h_sdram0_AWPROT  (f2h_sdram_slave_awprot),  //                 .awprot
		.f2h_sdram0_AWVALID (f2h_sdram_slave_awvalid), //                 .awvalid
		.f2h_sdram0_AWCACHE (f2h_sdram_slave_awcache), //                 .awcache
		.f2h_sdram0_BRESP   (f2h_sdram_slave_bresp),   //                 .bresp
		.f2h_sdram0_BID     (f2h_sdram_slave_bid),     //                 .bid
		.f2h_sdram0_BVALID  (f2h_sdram_slave_bvalid),  //                 .bvalid
		.f2h_sdram0_BREADY  (f2h_sdram_slave_bready),  //                 .bready
		.f2h_sdram0_ARREADY (f2h_sdram_slave_arready), //                 .arready
		.f2h_sdram0_AWREADY (f2h_sdram_slave_awready), //                 .awready
		.f2h_sdram0_RREADY  (f2h_sdram_slave_rready),  //                 .rready
		.f2h_sdram0_RDATA   (f2h_sdram_slave_rdata),   //                 .rdata
		.f2h_sdram0_RRESP   (f2h_sdram_slave_rresp),   //                 .rresp
		.f2h_sdram0_RLAST   (f2h_sdram_slave_rlast),   //                 .rlast
		.f2h_sdram0_RID     (f2h_sdram_slave_rid),     //                 .rid
		.f2h_sdram0_RVALID  (f2h_sdram_slave_rvalid),  //                 .rvalid
		.f2h_sdram0_WLAST   (f2h_sdram_slave_wlast),   //                 .wlast
		.f2h_sdram0_WVALID  (f2h_sdram_slave_wvalid),  //                 .wvalid
		.f2h_sdram0_WDATA   (f2h_sdram_slave_wdata),   //                 .wdata
		.f2h_sdram0_WSTRB   (f2h_sdram_slave_wstrb),   //                 .wstrb
		.f2h_sdram0_WREADY  (f2h_sdram_slave_wready),  //                 .wready
		.f2h_sdram0_WID     (f2h_sdram_slave_wid),     //                 .wid
		.h2f_axi_clk        (h2f_axi_clk_clk),         //    h2f_axi_clock.clk
		.h2f_AWID           (h2f_axi_master_awid),     //   h2f_axi_master.awid
		.h2f_AWADDR         (h2f_axi_master_awaddr),   //                 .awaddr
		.h2f_AWLEN          (h2f_axi_master_awlen),    //                 .awlen
		.h2f_AWSIZE         (h2f_axi_master_awsize),   //                 .awsize
		.h2f_AWBURST        (h2f_axi_master_awburst),  //                 .awburst
		.h2f_AWLOCK         (h2f_axi_master_awlock),   //                 .awlock
		.h2f_AWCACHE        (h2f_axi_master_awcache),  //                 .awcache
		.h2f_AWPROT         (h2f_axi_master_awprot),   //                 .awprot
		.h2f_AWVALID        (h2f_axi_master_awvalid),  //                 .awvalid
		.h2f_AWREADY        (h2f_axi_master_awready),  //                 .awready
		.h2f_WID            (h2f_axi_master_wid),      //                 .wid
		.h2f_WDATA          (h2f_axi_master_wdata),    //                 .wdata
		.h2f_WSTRB          (h2f_axi_master_wstrb),    //                 .wstrb
		.h2f_WLAST          (h2f_axi_master_wlast),    //                 .wlast
		.h2f_WVALID         (h2f_axi_master_wvalid),   //                 .wvalid
		.h2f_WREADY         (h2f_axi_master_wready),   //                 .wready
		.h2f_BID            (h2f_axi_master_bid),      //                 .bid
		.h2f_BRESP          (h2f_axi_master_bresp),    //                 .bresp
		.h2f_BVALID         (h2f_axi_master_bvalid),   //                 .bvalid
		.h2f_BREADY         (h2f_axi_master_bready),   //                 .bready
		.h2f_ARID           (h2f_axi_master_arid),     //                 .arid
		.h2f_ARADDR         (h2f_axi_master_araddr),   //                 .araddr
		.h2f_ARLEN          (h2f_axi_master_arlen),    //                 .arlen
		.h2f_ARSIZE         (h2f_axi_master_arsize),   //                 .arsize
		.h2f_ARBURST        (h2f_axi_master_arburst),  //                 .arburst
		.h2f_ARLOCK         (h2f_axi_master_arlock),   //                 .arlock
		.h2f_ARCACHE        (h2f_axi_master_arcache),  //                 .arcache
		.h2f_ARPROT         (h2f_axi_master_arprot),   //                 .arprot
		.h2f_ARVALID        (h2f_axi_master_arvalid),  //                 .arvalid
		.h2f_ARREADY        (h2f_axi_master_arready),  //                 .arready
		.h2f_RID            (h2f_axi_master_rid),      //                 .rid
		.h2f_RDATA          (h2f_axi_master_rdata),    //                 .rdata
		.h2f_RRESP          (h2f_axi_master_rresp),    //                 .rresp
		.h2f_RLAST          (h2f_axi_master_rlast),    //                 .rlast
		.h2f_RVALID         (h2f_axi_master_rvalid),   //                 .rvalid
		.h2f_RREADY         (h2f_axi_master_rready),   //                 .rready
		.f2h_irq_p0         (irq0_irq),                //         f2h_irq0.irq
		.f2h_irq_p1         (irq1_irq)                 //         f2h_irq1.irq
	);

endmodule
